module main

@[export: "square"]
fn square(i int) int {
	return i * i
}
